class OutData;
	bit sof;
	int llr_data;
	int extr_data;
	bit eof;
endclass