class Test6144 extends BaseTest;

	function new();
		ref_extrinsic_path = "./extrinsic_6144.txt";
		ref_llr_path       = "./LLR_6144.txt";
		stimuli_path       = "./in_6144.txt";
		test_name          = "6144";
	endfunction

endclass