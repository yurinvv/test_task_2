package tb_pckg;
	`include "Driver.svh"
	`include "OutData.svh"
	`include "Monitor.svh"
	`include "Scoreboard.svh"
	`include "Environment.svh"
	`include "BaseTest.svh"
	`include "Test512.svh"
	`include "Test6144.svh"
endpackage